magic
tech sky130A
magscale 1 2
timestamp 1611863236
<< nwell >>
rect 34003 -10491 34535 -9850
<< locali >>
rect 33817 -10573 33832 -10539
rect 33866 -10573 34131 -10539
rect 34449 -10584 35003 -10550
rect 35041 -10584 35057 -10550
rect 33972 -10890 34056 -10870
rect 33972 -10940 33993 -10890
rect 34035 -10940 34056 -10890
rect 33972 -10954 34056 -10940
rect 34554 -10885 34672 -10884
rect 34554 -10920 34625 -10885
rect 34659 -10920 34672 -10885
rect 34554 -10952 34574 -10920
<< viali >>
rect 34272 -10507 34310 -10471
rect 33832 -10573 33866 -10539
rect 35003 -10584 35041 -10550
rect 33993 -10940 34035 -10890
rect 34625 -10920 34659 -10885
<< metal1 >>
rect 34056 -9552 34142 -9542
rect 34056 -9626 34080 -9552
rect 34056 -9638 34142 -9626
rect 33875 -10144 34498 -10082
rect 33875 -10262 33910 -10144
rect 33968 -10262 34498 -10144
rect 33875 -10288 34498 -10262
rect 33875 -10289 34086 -10288
rect 34716 -10454 34780 -10448
rect 34249 -10465 34358 -10462
rect 34716 -10465 34722 -10454
rect 34249 -10471 34722 -10465
rect 34249 -10507 34272 -10471
rect 34310 -10506 34722 -10471
rect 34774 -10506 34780 -10454
rect 34310 -10507 34780 -10506
rect 34249 -10513 34780 -10507
rect 34716 -10514 34780 -10513
rect 33820 -10522 33890 -10516
rect 33820 -10574 33832 -10522
rect 33884 -10574 33890 -10522
rect 33820 -10584 33890 -10574
rect 34990 -10528 35070 -10516
rect 34990 -10550 35011 -10528
rect 34990 -10584 35003 -10550
rect 35064 -10580 35070 -10528
rect 35041 -10584 35070 -10580
rect 34990 -10596 35070 -10584
rect 34618 -10868 34684 -10862
rect 33972 -10888 34056 -10870
rect 33972 -10947 33986 -10888
rect 34044 -10947 34056 -10888
rect 34618 -10920 34625 -10868
rect 34678 -10920 34684 -10868
rect 34618 -10932 34684 -10920
rect 33972 -10954 34056 -10947
<< via1 >>
rect 34080 -9626 34160 -9552
rect 33910 -10262 33968 -10144
rect 34722 -10506 34774 -10454
rect 33832 -10539 33884 -10522
rect 33832 -10573 33866 -10539
rect 33866 -10573 33884 -10539
rect 33832 -10574 33884 -10573
rect 35011 -10550 35064 -10528
rect 35011 -10580 35041 -10550
rect 35041 -10580 35064 -10550
rect 33986 -10947 34044 -10888
rect 34625 -10885 34678 -10868
rect 34625 -10920 34659 -10885
rect 34659 -10920 34678 -10885
<< metal2 >>
rect 34056 -9542 34198 -9534
rect 34056 -9629 34073 -9542
rect 34186 -9629 34198 -9542
rect 34056 -9638 34198 -9629
rect 33875 -10126 34002 -10082
rect 33875 -10263 33908 -10126
rect 33970 -10263 34002 -10126
rect 33875 -10290 34002 -10263
rect 34712 -10450 34788 -10440
rect 34712 -10506 34722 -10450
rect 34778 -10506 34788 -10450
rect 33820 -10518 33898 -10508
rect 34712 -10516 34788 -10506
rect 33820 -10574 33832 -10518
rect 33888 -10574 33898 -10518
rect 33820 -10584 33898 -10574
rect 34990 -10528 35070 -10516
rect 34990 -10586 35003 -10528
rect 35064 -10580 35070 -10528
rect 35059 -10586 35070 -10580
rect 34990 -10596 35070 -10586
rect 34756 -10862 34840 -10854
rect 34619 -10864 34840 -10862
rect 33850 -10875 34056 -10864
rect 33850 -10941 33864 -10875
rect 33928 -10888 34056 -10875
rect 33928 -10941 33986 -10888
rect 33850 -10947 33986 -10941
rect 34044 -10947 34056 -10888
rect 34619 -10868 34762 -10864
rect 34619 -10920 34625 -10868
rect 34678 -10920 34762 -10868
rect 34619 -10922 34762 -10920
rect 34830 -10922 34840 -10864
rect 34619 -10926 34840 -10922
rect 33850 -10956 34056 -10947
<< via2 >>
rect 34073 -9552 34186 -9542
rect 34073 -9626 34080 -9552
rect 34080 -9626 34160 -9552
rect 34160 -9626 34186 -9552
rect 34073 -9629 34186 -9626
rect 33908 -10144 33970 -10126
rect 33908 -10262 33910 -10144
rect 33910 -10262 33968 -10144
rect 33968 -10262 33970 -10144
rect 33908 -10263 33970 -10262
rect 34722 -10454 34778 -10450
rect 34722 -10506 34774 -10454
rect 34774 -10506 34778 -10454
rect 33832 -10522 33888 -10518
rect 33832 -10574 33884 -10522
rect 33884 -10574 33888 -10522
rect 35003 -10580 35011 -10528
rect 35011 -10580 35059 -10528
rect 35003 -10586 35059 -10580
rect 33864 -10941 33928 -10875
rect 34762 -10922 34830 -10864
<< metal3 >>
rect 5345 -8213 20015 -8047
rect 5345 -22654 5511 -8213
rect 19042 -8846 19127 -8836
rect 19042 -8911 19058 -8846
rect 19122 -8911 19127 -8846
rect 19042 -10513 19127 -8911
rect 19849 -9502 20015 -8213
rect 19849 -9534 34089 -9502
rect 19849 -9542 34200 -9534
rect 19849 -9629 34073 -9542
rect 34186 -9629 34200 -9542
rect 19849 -9638 34200 -9629
rect 19849 -9668 34089 -9638
rect 33874 -10126 34002 -10082
rect 33874 -10264 33908 -10126
rect 33972 -10264 34002 -10126
rect 33874 -10290 34002 -10264
rect 34990 -10414 57135 -10392
rect 34713 -10428 34818 -10420
rect 34713 -10450 34741 -10428
rect 33747 -10513 33898 -10492
rect 19042 -10518 33898 -10513
rect 34713 -10506 34722 -10450
rect 34806 -10492 34818 -10428
rect 34778 -10506 34818 -10492
rect 34713 -10515 34818 -10506
rect 34990 -10486 57034 -10414
rect 57116 -10486 57135 -10414
rect 34990 -10498 57135 -10486
rect 19042 -10574 33832 -10518
rect 33888 -10574 33898 -10518
rect 19042 -10598 33898 -10574
rect 34990 -10528 35096 -10498
rect 34566 -10616 34642 -10584
rect 34990 -10586 35003 -10528
rect 35059 -10586 35096 -10528
rect 34990 -10598 35096 -10586
rect 34626 -10699 34642 -10616
rect 34566 -10734 34642 -10699
rect 33850 -10874 33940 -10842
rect 33850 -10942 33864 -10874
rect 33928 -10942 33940 -10874
rect 33850 -10956 33940 -10942
rect 34748 -10858 34852 -10826
rect 34748 -10864 34768 -10858
rect 34748 -10922 34762 -10864
rect 34748 -10924 34768 -10922
rect 34834 -10924 34852 -10858
rect 34748 -10950 34852 -10924
rect 34573 -11028 34592 -10968
rect 34580 -11092 34592 -11028
rect 34573 -11115 34592 -11092
rect 5345 -22756 5390 -22654
rect 5470 -22756 5511 -22654
rect 5345 -22783 5511 -22756
<< via3 >>
rect 19058 -8911 19122 -8846
rect 33908 -10263 33970 -10126
rect 33970 -10263 33972 -10126
rect 33908 -10264 33972 -10263
rect 34741 -10450 34806 -10428
rect 34741 -10492 34778 -10450
rect 34778 -10492 34806 -10450
rect 57034 -10486 57116 -10414
rect 34540 -10699 34626 -10616
rect 33864 -10875 33928 -10874
rect 33864 -10941 33928 -10875
rect 33864 -10942 33928 -10941
rect 34768 -10864 34834 -10858
rect 34768 -10922 34830 -10864
rect 34830 -10922 34834 -10864
rect 34768 -10924 34834 -10922
rect 34515 -11092 34580 -11028
rect 5390 -22756 5470 -22654
<< metal4 >>
rect 1811 -10092 2017 133
rect 19048 -8766 19128 52
rect 19044 -8846 19136 -8766
rect 19044 -8911 19058 -8846
rect 19122 -8911 19136 -8846
rect 19044 -8916 19136 -8911
rect 33761 -10092 34002 -10082
rect 1811 -10126 34002 -10092
rect 1811 -10264 33908 -10126
rect 33972 -10264 34002 -10126
rect 1811 -10290 34002 -10264
rect 1811 -10298 33937 -10290
rect 34726 -10318 34836 111
rect 34724 -10428 34836 -10318
rect 34724 -10492 34741 -10428
rect 34806 -10492 34836 -10428
rect 34724 -10514 34836 -10492
rect 34518 -10616 34700 -10584
rect 34518 -10699 34540 -10616
rect 34626 -10643 34700 -10616
rect 43741 -10643 43815 69
rect 57016 11 57485 133
rect 57016 -10414 57138 11
rect 57016 -10486 57034 -10414
rect 57116 -10486 57138 -10414
rect 57016 -10502 57138 -10486
rect 34626 -10699 43815 -10643
rect 34518 -10717 43815 -10699
rect 34518 -10734 34700 -10717
rect 33850 -10874 33940 -10842
rect 33850 -10942 33864 -10874
rect 33928 -10942 33940 -10874
rect 33850 -10966 33940 -10942
rect 33849 -10995 33940 -10966
rect 34758 -10858 34842 -10830
rect 34758 -10924 34768 -10858
rect 34834 -10924 34842 -10858
rect 33849 -17566 33913 -10995
rect 34506 -11028 34590 -11020
rect 34506 -11092 34515 -11028
rect 34580 -11092 34590 -11028
rect 34506 -11112 34590 -11092
rect 34506 -11216 34572 -11112
rect 24314 -17630 33913 -17566
rect 5345 -22654 5512 -22632
rect 5345 -22756 5390 -22654
rect 5470 -22756 5512 -22654
rect 5345 -22826 5512 -22756
rect 5345 -22883 5514 -22826
rect 5346 -24994 5514 -22883
rect 24314 -25006 24378 -17630
rect 34508 -24943 34570 -11216
rect 34758 -17488 34842 -10924
rect 34758 -17572 43404 -17488
rect 43320 -25008 43404 -17572
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_11 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1611854809
transform 1 0 540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_10
timestamp 1611854809
transform 1 0 14540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_9
timestamp 1611854809
transform 1 0 28540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_8
timestamp 1611854809
transform 1 0 42540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_7
timestamp 1611854809
transform 1 0 56540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_6
timestamp 1611854809
transform 1 0 70540 0 -1 -25460
box -540 -540 12540 14540
use BITCELL  BITCELL_0
timestamp 1611860754
transform 1 0 33491 0 1 -10948
box 515 -167 1083 753
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611854809
transform 1 0 34106 0 -1 -9590
box -38 -48 130 592
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_0
timestamp 1611854809
transform 1 0 540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_1
timestamp 1611854809
transform 1 0 14540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_3
timestamp 1611854809
transform 1 0 28540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_2
timestamp 1611854809
transform 1 0 42540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_5
timestamp 1611854809
transform 1 0 56540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_4
timestamp 1611854809
transform 1 0 70540 0 1 540
box -540 -540 12540 14540
<< labels >>
flabel space 384 390 384 390 1 FreeSans 6400 0 0 0 VDD
flabel space 14394 400 14394 400 1 FreeSans 6400 0 0 0 Q
flabel space 28406 392 28406 392 1 FreeSans 6400 0 0 0 SENSE_N
flabel space 42400 400 42400 400 1 FreeSans 6400 0 0 0 BLB
flabel space 56414 392 56414 392 1 FreeSans 6400 0 0 0 QN
flabel space 418 -39598 418 -39598 1 FreeSans 6400 0 0 0 VSS
flabel space 14406 -39596 14406 -39596 1 FreeSans 6400 0 0 0 WRR
flabel space 28410 -39596 28410 -39596 1 FreeSans 6400 0 0 0 BL
flabel space 42398 -39608 42398 -39608 1 FreeSans 6400 0 0 0 WRL
<< end >>
