magic
tech sky130A
magscale 1 2
timestamp 1612375005
<< nwell >>
rect 34004 -9850 35650 -9848
rect 34003 -10491 35650 -9850
rect 34004 -10492 35650 -10491
<< locali >>
rect 34272 -10472 34310 -10471
rect 34272 -10506 34274 -10472
rect 34308 -10506 34310 -10472
rect 34272 -10507 34310 -10506
rect 33665 -10573 33680 -10539
rect 33714 -10573 34131 -10539
rect 35172 -10548 35240 -10542
rect 34449 -10569 34514 -10550
rect 34449 -10584 34479 -10569
rect 34452 -10603 34479 -10584
rect 34513 -10584 34514 -10569
rect 35172 -10582 35188 -10548
rect 35222 -10582 35240 -10548
rect 35172 -10584 35240 -10582
rect 34513 -10603 34530 -10584
rect 35559 -10585 35639 -10551
rect 35673 -10585 35689 -10551
rect 34452 -10630 34530 -10603
rect 33972 -10898 34056 -10870
rect 33972 -10932 33997 -10898
rect 34031 -10932 34056 -10898
rect 33972 -10954 34056 -10932
rect 34554 -10886 34672 -10884
rect 34554 -10920 34625 -10886
rect 34659 -10920 34672 -10886
rect 35070 -10902 35166 -10886
rect 34554 -10952 34574 -10920
rect 35070 -10936 35080 -10902
rect 35114 -10936 35166 -10902
rect 35070 -10954 35166 -10936
rect 35634 -10901 35748 -10884
rect 35634 -10935 35699 -10901
rect 35733 -10935 35748 -10901
rect 35634 -10953 35748 -10935
<< viali >>
rect 34274 -10506 34308 -10472
rect 33680 -10573 33714 -10539
rect 34479 -10603 34513 -10569
rect 35188 -10582 35222 -10548
rect 35639 -10585 35673 -10551
rect 33997 -10932 34031 -10898
rect 34625 -10920 34659 -10886
rect 35080 -10936 35114 -10902
rect 35699 -10935 35733 -10901
<< metal1 >>
rect 34056 -9552 34142 -9542
rect 34056 -9563 34160 -9552
rect 34056 -9615 34094 -9563
rect 34146 -9615 34160 -9563
rect 34056 -9626 34160 -9615
rect 34056 -9638 34142 -9626
rect 33875 -10145 35775 -10082
rect 33875 -10197 33913 -10145
rect 33965 -10197 35775 -10145
rect 33875 -10209 35775 -10197
rect 33875 -10261 33913 -10209
rect 33965 -10261 35775 -10209
rect 33875 -10288 35775 -10261
rect 33875 -10289 34086 -10288
rect 34206 -10289 35775 -10288
rect 34716 -10454 34780 -10448
rect 34249 -10465 34358 -10462
rect 34716 -10465 34722 -10454
rect 34249 -10472 34722 -10465
rect 34249 -10506 34274 -10472
rect 34308 -10506 34722 -10472
rect 34774 -10465 34780 -10454
rect 34774 -10506 35452 -10465
rect 34249 -10513 35452 -10506
rect 34716 -10514 34780 -10513
rect 33668 -10522 33738 -10516
rect 33668 -10574 33680 -10522
rect 33732 -10574 33738 -10522
rect 35704 -10534 35768 -10528
rect 35704 -10536 35710 -10534
rect 35003 -10548 35234 -10542
rect 33668 -10584 33738 -10574
rect 34454 -10558 34532 -10550
rect 34454 -10610 34476 -10558
rect 34528 -10610 34532 -10558
rect 35003 -10584 35010 -10548
rect 35004 -10600 35010 -10584
rect 35062 -10582 35188 -10548
rect 35222 -10582 35234 -10548
rect 35062 -10590 35234 -10582
rect 35624 -10551 35710 -10536
rect 35624 -10585 35639 -10551
rect 35673 -10585 35710 -10551
rect 35624 -10586 35710 -10585
rect 35762 -10586 35768 -10534
rect 35062 -10600 35068 -10590
rect 35624 -10594 35768 -10586
rect 35004 -10606 35068 -10600
rect 34454 -10628 34532 -10610
rect 34618 -10868 34684 -10862
rect 33972 -10892 34056 -10870
rect 33972 -10944 33989 -10892
rect 34041 -10944 34056 -10892
rect 34618 -10920 34625 -10868
rect 34677 -10920 34684 -10868
rect 34618 -10932 34684 -10920
rect 35012 -10892 35130 -10886
rect 33972 -10954 34056 -10944
rect 35012 -10944 35019 -10892
rect 35071 -10902 35130 -10892
rect 35071 -10936 35080 -10902
rect 35114 -10936 35130 -10902
rect 35071 -10944 35130 -10936
rect 35012 -10954 35130 -10944
rect 35682 -10893 35852 -10884
rect 35682 -10901 35776 -10893
rect 35682 -10935 35699 -10901
rect 35733 -10935 35776 -10901
rect 35682 -10945 35776 -10935
rect 35828 -10945 35852 -10893
rect 35682 -10952 35852 -10945
<< via1 >>
rect 34094 -9615 34146 -9563
rect 33913 -10197 33965 -10145
rect 33913 -10261 33965 -10209
rect 34722 -10506 34774 -10454
rect 33680 -10539 33732 -10522
rect 33680 -10573 33714 -10539
rect 33714 -10573 33732 -10539
rect 33680 -10574 33732 -10573
rect 34476 -10569 34528 -10558
rect 34476 -10603 34479 -10569
rect 34479 -10603 34513 -10569
rect 34513 -10603 34528 -10569
rect 34476 -10610 34528 -10603
rect 35010 -10600 35062 -10548
rect 35710 -10586 35762 -10534
rect 33989 -10898 34041 -10892
rect 33989 -10932 33997 -10898
rect 33997 -10932 34031 -10898
rect 34031 -10932 34041 -10898
rect 33989 -10944 34041 -10932
rect 34625 -10886 34677 -10868
rect 34625 -10920 34659 -10886
rect 34659 -10920 34677 -10886
rect 35019 -10944 35071 -10892
rect 35776 -10945 35828 -10893
<< metal2 >>
rect 34456 -9516 34586 -9504
rect 34056 -9558 34198 -9534
rect 34056 -9563 34101 -9558
rect 34056 -9615 34094 -9563
rect 34157 -9614 34198 -9558
rect 34456 -9572 34503 -9516
rect 34559 -9572 34586 -9516
rect 34456 -9608 34586 -9572
rect 34146 -9615 34198 -9614
rect 34056 -9638 34198 -9615
rect 33875 -10127 34002 -10082
rect 33875 -10183 33911 -10127
rect 33967 -10183 34002 -10127
rect 33875 -10197 33913 -10183
rect 33965 -10197 34002 -10183
rect 33875 -10207 34002 -10197
rect 33875 -10263 33911 -10207
rect 33967 -10263 34002 -10207
rect 33875 -10290 34002 -10263
rect 33668 -10518 33746 -10508
rect 33668 -10574 33680 -10518
rect 33736 -10574 33746 -10518
rect 34464 -10550 34504 -9608
rect 34984 -9708 35064 -9700
rect 34984 -9764 34994 -9708
rect 35050 -9764 35064 -9708
rect 34984 -9772 35064 -9764
rect 34712 -10450 34788 -10440
rect 34712 -10506 34722 -10450
rect 34778 -10506 34788 -10450
rect 34712 -10516 34788 -10506
rect 35004 -10542 35033 -9772
rect 35704 -9872 35802 -9846
rect 35704 -9928 35728 -9872
rect 35784 -9928 35802 -9872
rect 35704 -9952 35802 -9928
rect 35704 -10528 35764 -9952
rect 35704 -10534 35768 -10528
rect 35004 -10548 35068 -10542
rect 33668 -10584 33746 -10574
rect 34456 -10558 34532 -10550
rect 34456 -10610 34476 -10558
rect 34528 -10610 34532 -10558
rect 35004 -10600 35010 -10548
rect 35062 -10600 35068 -10548
rect 35704 -10586 35710 -10534
rect 35762 -10586 35768 -10534
rect 35704 -10592 35768 -10586
rect 35004 -10606 35068 -10600
rect 34456 -10630 34532 -10610
rect 33850 -10880 34056 -10864
rect 33850 -10936 33868 -10880
rect 33924 -10892 34056 -10880
rect 33924 -10936 33989 -10892
rect 33850 -10944 33989 -10936
rect 34041 -10944 34056 -10892
rect 34619 -10868 34678 -10862
rect 34619 -10920 34625 -10868
rect 34677 -10920 34678 -10868
rect 35770 -10883 35956 -10874
rect 34619 -10926 34678 -10920
rect 35012 -10892 35078 -10886
rect 33850 -10956 34056 -10944
rect 34624 -11342 34664 -10926
rect 35012 -10944 35019 -10892
rect 35071 -10944 35078 -10892
rect 35012 -10954 35078 -10944
rect 35770 -10893 35883 -10883
rect 35770 -10945 35776 -10893
rect 35828 -10939 35883 -10893
rect 35939 -10939 35956 -10883
rect 35828 -10945 35956 -10939
rect 35770 -10954 35956 -10945
rect 35018 -10962 35070 -10954
rect 35024 -11232 35057 -10962
rect 35024 -11233 35096 -11232
rect 35021 -11238 35097 -11233
rect 35021 -11294 35030 -11238
rect 35086 -11294 35097 -11238
rect 35021 -11303 35097 -11294
rect 34732 -11342 34880 -11316
rect 34624 -11350 34880 -11342
rect 34624 -11406 34774 -11350
rect 34830 -11406 34880 -11350
rect 34624 -11422 34880 -11406
rect 34732 -11452 34880 -11422
<< via2 >>
rect 34101 -9563 34157 -9558
rect 34101 -9614 34146 -9563
rect 34146 -9614 34157 -9563
rect 34503 -9572 34559 -9516
rect 33911 -10145 33967 -10127
rect 33911 -10183 33913 -10145
rect 33913 -10183 33965 -10145
rect 33965 -10183 33967 -10145
rect 33911 -10209 33967 -10207
rect 33911 -10261 33913 -10209
rect 33913 -10261 33965 -10209
rect 33965 -10261 33967 -10209
rect 33911 -10263 33967 -10261
rect 33680 -10522 33736 -10518
rect 33680 -10574 33732 -10522
rect 33732 -10574 33736 -10522
rect 34994 -9764 35050 -9708
rect 34722 -10454 34778 -10450
rect 34722 -10506 34774 -10454
rect 34774 -10506 34778 -10454
rect 35728 -9928 35784 -9872
rect 33868 -10936 33924 -10880
rect 35883 -10939 35939 -10883
rect 35030 -11294 35086 -11238
rect 34774 -11406 34830 -11350
<< metal3 >>
rect 19849 -9502 20015 -9501
rect 5363 -9534 34089 -9502
rect 34446 -9506 34618 -9466
rect 56876 -9502 57168 -9488
rect 56866 -9506 57168 -9502
rect 34446 -9516 57168 -9506
rect 5363 -9556 34200 -9534
rect 5363 -9620 5419 -9556
rect 5483 -9558 34200 -9556
rect 5483 -9614 34101 -9558
rect 34157 -9614 34200 -9558
rect 5483 -9620 34200 -9614
rect 34446 -9572 34503 -9516
rect 34559 -9532 57168 -9516
rect 34559 -9572 57041 -9532
rect 34446 -9596 57041 -9572
rect 57105 -9596 57168 -9532
rect 34446 -9612 57168 -9596
rect 34446 -9618 34998 -9612
rect 56866 -9616 57168 -9612
rect 5363 -9638 34200 -9620
rect 56876 -9628 57168 -9616
rect 5363 -9668 34089 -9638
rect 74238 -9685 74370 -9670
rect 34984 -9701 35064 -9698
rect 74238 -9701 74283 -9685
rect 34984 -9708 74283 -9701
rect 34984 -9764 34994 -9708
rect 35050 -9749 74283 -9708
rect 74347 -9749 74370 -9685
rect 35050 -9764 74370 -9749
rect 34984 -9767 74370 -9764
rect 34984 -9770 35064 -9767
rect 74238 -9796 74370 -9767
rect 35708 -9866 87016 -9864
rect 35708 -9872 87137 -9866
rect 35708 -9928 35728 -9872
rect 35784 -9928 87137 -9872
rect 35708 -9930 87137 -9928
rect 87201 -9930 87300 -9866
rect 35708 -9938 87300 -9930
rect 35708 -9940 86968 -9938
rect 1764 -10053 4706 -10050
rect 17896 -10052 33980 -10050
rect 17896 -10053 34046 -10052
rect 1764 -10117 34046 -10053
rect 1764 -10261 1830 -10117
rect 2214 -10127 34046 -10117
rect 2214 -10183 33911 -10127
rect 33967 -10183 34046 -10127
rect 2214 -10207 34046 -10183
rect 2214 -10261 33911 -10207
rect 1764 -10263 33911 -10261
rect 33967 -10263 34046 -10207
rect 1764 -10318 34046 -10263
rect 33784 -10320 34046 -10318
rect 34713 -10428 34818 -10420
rect 34713 -10450 34741 -10428
rect 19042 -10513 19127 -10512
rect 33595 -10513 33746 -10492
rect 19042 -10518 33746 -10513
rect 34713 -10506 34722 -10450
rect 34805 -10492 34818 -10428
rect 34778 -10506 34818 -10492
rect 34713 -10515 34818 -10506
rect 19042 -10524 33680 -10518
rect 19042 -10588 19056 -10524
rect 19120 -10574 33680 -10524
rect 33736 -10574 33746 -10518
rect 19120 -10588 33746 -10574
rect 19042 -10598 33746 -10588
rect 34530 -10622 43859 -10586
rect 34530 -10686 43714 -10622
rect 43778 -10686 43859 -10622
rect 34530 -10732 43859 -10686
rect 33850 -10876 33940 -10842
rect 33850 -10940 33864 -10876
rect 33928 -10940 33940 -10876
rect 33850 -10956 33940 -10940
rect 35864 -10880 74600 -10870
rect 35864 -10883 74470 -10880
rect 35864 -10939 35883 -10883
rect 35939 -10939 74470 -10883
rect 35864 -10944 74470 -10939
rect 74534 -10944 74600 -10880
rect 35864 -10955 74600 -10944
rect 34506 -11114 35694 -10968
rect 34506 -11116 34624 -11114
rect 34506 -11184 34598 -11116
rect 34506 -11248 34516 -11184
rect 34580 -11248 34598 -11184
rect 59740 -11215 59922 -11168
rect 59740 -11232 59804 -11215
rect 34506 -11264 34598 -11248
rect 35022 -11238 59804 -11232
rect 35022 -11294 35030 -11238
rect 35086 -11279 59804 -11238
rect 59868 -11279 59922 -11215
rect 35086 -11294 59922 -11279
rect 35022 -11300 59922 -11294
rect 35022 -11302 35102 -11300
rect 34730 -11346 34878 -11316
rect 59740 -11328 59922 -11300
rect 34730 -11410 34770 -11346
rect 34834 -11410 34878 -11346
rect 34730 -11452 34878 -11410
<< via3 >>
rect 5419 -9620 5483 -9556
rect 57041 -9596 57105 -9532
rect 74283 -9749 74347 -9685
rect 87137 -9930 87201 -9866
rect 1830 -10261 2214 -10117
rect 34741 -10450 34805 -10428
rect 34741 -10492 34778 -10450
rect 34778 -10492 34805 -10450
rect 19056 -10588 19120 -10524
rect 43714 -10686 43778 -10622
rect 33864 -10880 33928 -10876
rect 33864 -10936 33868 -10880
rect 33868 -10936 33924 -10880
rect 33924 -10936 33928 -10880
rect 33864 -10940 33928 -10936
rect 74470 -10944 74534 -10880
rect 34516 -11248 34580 -11184
rect 59804 -11279 59868 -11215
rect 34770 -11350 34834 -11346
rect 34770 -11406 34774 -11350
rect 34774 -11406 34830 -11350
rect 34830 -11406 34834 -11350
rect 34770 -11410 34834 -11406
<< metal4 >>
rect 1811 -9792 2017 133
rect 19048 -8601 19128 52
rect 5363 -9556 5550 -9500
rect 5363 -9620 5419 -9556
rect 5483 -9620 5550 -9556
rect 1762 -10117 2288 -9792
rect 1762 -10261 1830 -10117
rect 2214 -10261 2288 -10117
rect 1762 -10320 2288 -10261
rect 5363 -23086 5550 -9620
rect 19040 -10524 19130 -8601
rect 34726 -10318 34836 111
rect 34724 -10428 34836 -10318
rect 34724 -10492 34741 -10428
rect 34805 -10492 34836 -10428
rect 34724 -10514 34836 -10492
rect 19040 -10588 19056 -10524
rect 19120 -10588 19130 -10524
rect 43665 -10538 43819 99
rect 57016 11 57485 133
rect 57016 -9400 57138 11
rect 74248 -150 74398 452
rect 56994 -9462 57188 -9400
rect 56992 -9532 57188 -9462
rect 56992 -9596 57041 -9532
rect 57105 -9596 57188 -9532
rect 74280 -9556 74352 -150
rect 56992 -9644 57188 -9596
rect 56994 -9650 57188 -9644
rect 74202 -9685 74432 -9556
rect 74202 -9749 74283 -9685
rect 74347 -9749 74432 -9685
rect 74202 -9816 74432 -9749
rect 87071 -9854 87301 477
rect 87071 -9866 87300 -9854
rect 87071 -9930 87137 -9866
rect 87201 -9930 87300 -9866
rect 87071 -9938 87300 -9930
rect 19040 -10602 19130 -10588
rect 43652 -10622 43854 -10538
rect 43652 -10686 43714 -10622
rect 43778 -10686 43854 -10622
rect 43652 -10734 43854 -10686
rect 33850 -10876 33940 -10842
rect 33850 -10940 33864 -10876
rect 33928 -10940 33940 -10876
rect 33850 -10966 33940 -10940
rect 74424 -10880 74600 -10870
rect 74424 -10944 74470 -10880
rect 74534 -10944 74600 -10880
rect 74424 -10955 74600 -10944
rect 74474 -10966 74544 -10955
rect 33849 -10995 33940 -10966
rect 33849 -17566 33913 -10995
rect 5346 -23274 5550 -23086
rect 24314 -17630 33913 -17566
rect 34500 -11184 34598 -11156
rect 34500 -11248 34516 -11184
rect 34580 -11248 34598 -11184
rect 5346 -24994 5514 -23274
rect 24314 -25006 24378 -17630
rect 34500 -24943 34598 -11248
rect 59740 -11215 59926 -11186
rect 59740 -11279 59804 -11215
rect 59868 -11279 59926 -11215
rect 34732 -11346 34878 -11316
rect 59740 -11328 59926 -11279
rect 34732 -11410 34770 -11346
rect 34834 -11410 34878 -11346
rect 34732 -11452 34878 -11410
rect 34758 -17488 34842 -11452
rect 34758 -17572 43404 -17488
rect 43320 -25008 43404 -17572
rect 59795 -25033 59861 -11328
rect 74477 -25503 74544 -10966
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_13
timestamp 1612207292
transform 1 0 540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_12
timestamp 1612207292
transform 1 0 14540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_11
timestamp 1612207292
transform 1 0 28540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_10
timestamp 1612207292
transform 1 0 42540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_9
timestamp 1612207292
transform 1 0 56540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_8
timestamp 1612207292
transform 1 0 70540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_7
timestamp 1612207292
transform 1 0 84540 0 -1 -25460
box -540 -540 12540 14540
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0
timestamp 1612207292
transform 1 0 34106 0 -1 -9590
box -38 -48 130 592
use BITCELL  BITCELL_0
timestamp 1612374967
transform 1 0 33491 0 1 -10948
box 515 -167 1083 753
use BITCELL  BITCELL_1
timestamp 1612374967
transform 1 0 34601 0 1 -10949
box 515 -167 1083 753
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_6
timestamp 1612207292
transform 1 0 540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_5
timestamp 1612207292
transform 1 0 14540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_4
timestamp 1612207292
transform 1 0 28540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_3
timestamp 1612207292
transform 1 0 42540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_2
timestamp 1612207292
transform 1 0 56540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_1
timestamp 1612207292
transform 1 0 70540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_0
timestamp 1612207292
transform 1 0 84540 0 1 540
box -540 -540 12540 14540
<< end >>
