magic
tech sky130A
magscale 1 2
timestamp 1611950381
<< nwell >>
rect 34004 -9850 35650 -9848
rect 34003 -10491 35650 -9850
rect 34004 -10492 35650 -10491
<< locali >>
rect 33665 -10573 33680 -10539
rect 33714 -10573 34131 -10539
rect 35172 -10548 35240 -10542
rect 34449 -10566 34514 -10550
rect 34449 -10584 34478 -10566
rect 34452 -10606 34478 -10584
rect 35172 -10582 35188 -10548
rect 35222 -10582 35240 -10548
rect 35172 -10584 35240 -10582
rect 34514 -10606 34530 -10584
rect 35559 -10585 35639 -10551
rect 35673 -10585 35689 -10551
rect 34452 -10630 34530 -10606
rect 33972 -10890 34056 -10870
rect 33972 -10940 33993 -10890
rect 34035 -10940 34056 -10890
rect 33972 -10954 34056 -10940
rect 34554 -10885 34672 -10884
rect 34554 -10920 34625 -10885
rect 34659 -10920 34672 -10885
rect 35070 -10902 35166 -10886
rect 34554 -10952 34574 -10920
rect 35070 -10936 35080 -10902
rect 35114 -10936 35166 -10902
rect 35070 -10954 35166 -10936
rect 35634 -10898 35748 -10884
rect 35634 -10938 35696 -10898
rect 35736 -10938 35748 -10898
rect 35634 -10953 35748 -10938
<< viali >>
rect 34272 -10507 34310 -10471
rect 33680 -10573 33714 -10539
rect 34478 -10606 34514 -10566
rect 35188 -10582 35222 -10548
rect 35639 -10585 35673 -10551
rect 33993 -10940 34035 -10890
rect 34625 -10920 34659 -10885
rect 35080 -10936 35114 -10902
rect 35696 -10938 35736 -10898
<< metal1 >>
rect 34056 -9552 34142 -9542
rect 34056 -9626 34080 -9552
rect 34056 -9638 34142 -9626
rect 33875 -10144 35775 -10082
rect 33875 -10262 33910 -10144
rect 33968 -10262 35775 -10144
rect 33875 -10288 35775 -10262
rect 33875 -10289 34086 -10288
rect 34206 -10289 35775 -10288
rect 34716 -10454 34780 -10448
rect 34249 -10465 34358 -10462
rect 34716 -10465 34722 -10454
rect 34249 -10471 34722 -10465
rect 34249 -10507 34272 -10471
rect 34310 -10506 34722 -10471
rect 34774 -10465 34780 -10454
rect 34774 -10506 35452 -10465
rect 34310 -10507 35452 -10506
rect 34249 -10513 35452 -10507
rect 34716 -10514 34780 -10513
rect 33668 -10522 33738 -10516
rect 33668 -10574 33680 -10522
rect 33732 -10574 33738 -10522
rect 35704 -10534 35768 -10528
rect 35704 -10536 35710 -10534
rect 35003 -10548 35234 -10542
rect 33668 -10584 33738 -10574
rect 34454 -10558 34532 -10550
rect 34454 -10610 34476 -10558
rect 34528 -10610 34532 -10558
rect 35003 -10584 35010 -10548
rect 35004 -10600 35010 -10584
rect 35062 -10582 35188 -10548
rect 35222 -10582 35234 -10548
rect 35062 -10590 35234 -10582
rect 35624 -10551 35710 -10536
rect 35624 -10585 35639 -10551
rect 35673 -10585 35710 -10551
rect 35624 -10586 35710 -10585
rect 35762 -10586 35768 -10534
rect 35062 -10600 35068 -10590
rect 35624 -10594 35768 -10586
rect 35004 -10606 35068 -10600
rect 34454 -10628 34532 -10610
rect 34618 -10868 34684 -10862
rect 33972 -10888 34056 -10870
rect 33972 -10947 33986 -10888
rect 34044 -10947 34056 -10888
rect 34618 -10920 34625 -10868
rect 34678 -10920 34684 -10868
rect 34618 -10932 34684 -10920
rect 35012 -10892 35130 -10886
rect 33972 -10954 34056 -10947
rect 35012 -10944 35019 -10892
rect 35071 -10902 35130 -10892
rect 35071 -10936 35080 -10902
rect 35114 -10936 35130 -10902
rect 35071 -10944 35130 -10936
rect 35012 -10954 35130 -10944
rect 35682 -10893 35852 -10884
rect 35682 -10898 35776 -10893
rect 35682 -10938 35696 -10898
rect 35736 -10938 35776 -10898
rect 35682 -10945 35776 -10938
rect 35828 -10945 35852 -10893
rect 35682 -10952 35852 -10945
<< via1 >>
rect 34080 -9626 34160 -9552
rect 33910 -10262 33968 -10144
rect 34722 -10506 34774 -10454
rect 33680 -10539 33732 -10522
rect 33680 -10573 33714 -10539
rect 33714 -10573 33732 -10539
rect 33680 -10574 33732 -10573
rect 34476 -10566 34528 -10558
rect 34476 -10606 34478 -10566
rect 34478 -10606 34514 -10566
rect 34514 -10606 34528 -10566
rect 34476 -10610 34528 -10606
rect 35010 -10600 35062 -10548
rect 35710 -10586 35762 -10534
rect 33986 -10890 34044 -10888
rect 33986 -10940 33993 -10890
rect 33993 -10940 34035 -10890
rect 34035 -10940 34044 -10890
rect 33986 -10947 34044 -10940
rect 34625 -10885 34678 -10868
rect 34625 -10920 34659 -10885
rect 34659 -10920 34678 -10885
rect 35019 -10944 35071 -10892
rect 35776 -10945 35828 -10893
<< metal2 >>
rect 34456 -9516 34586 -9504
rect 34056 -9542 34198 -9534
rect 34056 -9629 34073 -9542
rect 34186 -9629 34198 -9542
rect 34456 -9572 34496 -9516
rect 34566 -9572 34586 -9516
rect 34456 -9608 34586 -9572
rect 34056 -9638 34198 -9629
rect 33875 -10126 34002 -10082
rect 33875 -10263 33908 -10126
rect 33970 -10263 34002 -10126
rect 33875 -10290 34002 -10263
rect 33668 -10518 33746 -10508
rect 33668 -10574 33680 -10518
rect 33736 -10574 33746 -10518
rect 34464 -10550 34504 -9608
rect 34984 -9708 35064 -9700
rect 34984 -9764 34994 -9708
rect 35050 -9764 35064 -9708
rect 34984 -9772 35064 -9764
rect 34712 -10450 34788 -10440
rect 34712 -10506 34722 -10450
rect 34778 -10506 34788 -10450
rect 34712 -10516 34788 -10506
rect 35004 -10542 35033 -9772
rect 35704 -9872 35802 -9846
rect 35704 -9928 35728 -9872
rect 35784 -9928 35802 -9872
rect 35704 -9952 35802 -9928
rect 35704 -10528 35764 -9952
rect 35704 -10534 35768 -10528
rect 35004 -10548 35068 -10542
rect 33668 -10584 33746 -10574
rect 34456 -10558 34532 -10550
rect 34456 -10610 34476 -10558
rect 34528 -10610 34532 -10558
rect 35004 -10600 35010 -10548
rect 35062 -10600 35068 -10548
rect 35704 -10586 35710 -10534
rect 35762 -10586 35768 -10534
rect 35704 -10592 35768 -10586
rect 35004 -10606 35068 -10600
rect 34456 -10630 34532 -10610
rect 33850 -10875 34056 -10864
rect 33850 -10941 33864 -10875
rect 33928 -10888 34056 -10875
rect 33928 -10941 33986 -10888
rect 33850 -10947 33986 -10941
rect 34044 -10947 34056 -10888
rect 34619 -10868 34678 -10862
rect 34619 -10920 34625 -10868
rect 35770 -10880 35956 -10874
rect 34619 -10926 34678 -10920
rect 35012 -10892 35078 -10886
rect 33850 -10956 34056 -10947
rect 34624 -11342 34664 -10926
rect 35012 -10944 35019 -10892
rect 35071 -10944 35078 -10892
rect 35012 -10954 35078 -10944
rect 35770 -10893 35876 -10880
rect 35770 -10945 35776 -10893
rect 35828 -10942 35876 -10893
rect 35946 -10942 35956 -10880
rect 35828 -10945 35956 -10942
rect 35770 -10954 35956 -10945
rect 35018 -10962 35070 -10954
rect 35024 -11232 35057 -10962
rect 35024 -11233 35096 -11232
rect 35021 -11238 35097 -11233
rect 35021 -11294 35030 -11238
rect 35086 -11294 35097 -11238
rect 35021 -11303 35097 -11294
rect 34732 -11342 34880 -11316
rect 34624 -11344 34880 -11342
rect 34624 -11412 34768 -11344
rect 34836 -11412 34880 -11344
rect 34624 -11422 34880 -11412
rect 34732 -11452 34880 -11422
<< via2 >>
rect 34073 -9552 34186 -9542
rect 34073 -9626 34080 -9552
rect 34080 -9626 34160 -9552
rect 34160 -9626 34186 -9552
rect 34073 -9629 34186 -9626
rect 34496 -9572 34566 -9516
rect 33908 -10144 33970 -10126
rect 33908 -10262 33910 -10144
rect 33910 -10262 33968 -10144
rect 33968 -10262 33970 -10144
rect 33908 -10263 33970 -10262
rect 33680 -10522 33736 -10518
rect 33680 -10574 33732 -10522
rect 33732 -10574 33736 -10522
rect 34994 -9764 35050 -9708
rect 34722 -10454 34778 -10450
rect 34722 -10506 34774 -10454
rect 34774 -10506 34778 -10454
rect 35728 -9928 35784 -9872
rect 33864 -10941 33928 -10875
rect 35876 -10942 35946 -10880
rect 35030 -11294 35086 -11238
rect 34768 -11412 34836 -11344
<< metal3 >>
rect 19849 -9502 20015 -9501
rect 5363 -9522 34089 -9502
rect 5363 -9654 5384 -9522
rect 5518 -9534 34089 -9522
rect 34446 -9506 34618 -9466
rect 56876 -9502 57168 -9488
rect 56866 -9506 57168 -9502
rect 34446 -9516 57168 -9506
rect 5518 -9542 34200 -9534
rect 5518 -9629 34073 -9542
rect 34186 -9629 34200 -9542
rect 34446 -9572 34496 -9516
rect 34566 -9528 57168 -9516
rect 34566 -9572 57032 -9528
rect 34446 -9600 57032 -9572
rect 57114 -9600 57168 -9528
rect 34446 -9612 57168 -9600
rect 34446 -9618 34998 -9612
rect 56866 -9616 57168 -9612
rect 56876 -9628 57168 -9616
rect 5518 -9638 34200 -9629
rect 5518 -9654 34089 -9638
rect 5363 -9668 34089 -9654
rect 74238 -9684 74370 -9670
rect 34984 -9701 35064 -9698
rect 74238 -9701 74282 -9684
rect 34984 -9708 74282 -9701
rect 34984 -9764 34994 -9708
rect 35050 -9750 74282 -9708
rect 74348 -9750 74370 -9684
rect 35050 -9764 74370 -9750
rect 34984 -9767 74370 -9764
rect 34984 -9770 35064 -9767
rect 74238 -9796 74370 -9767
rect 35708 -9866 87016 -9864
rect 35708 -9872 87118 -9866
rect 35708 -9928 35728 -9872
rect 35784 -9928 87118 -9872
rect 35708 -9930 87118 -9928
rect 87220 -9930 87300 -9866
rect 35708 -9938 87300 -9930
rect 35708 -9940 86968 -9938
rect 1764 -10053 4706 -10050
rect 17896 -10052 33980 -10050
rect 17896 -10053 34046 -10052
rect 1764 -10092 34046 -10053
rect 1764 -10286 1814 -10092
rect 2230 -10126 34046 -10092
rect 2230 -10263 33908 -10126
rect 33970 -10263 34046 -10126
rect 2230 -10286 34046 -10263
rect 1764 -10318 34046 -10286
rect 33784 -10320 34046 -10318
rect 34713 -10428 34818 -10420
rect 34713 -10450 34741 -10428
rect 19042 -10513 19127 -10512
rect 33595 -10513 33746 -10492
rect 19042 -10518 33746 -10513
rect 34713 -10506 34722 -10450
rect 34806 -10492 34818 -10428
rect 34778 -10506 34818 -10492
rect 34713 -10515 34818 -10506
rect 19042 -10524 33680 -10518
rect 19042 -10588 19056 -10524
rect 19120 -10574 33680 -10524
rect 33736 -10574 33746 -10518
rect 19120 -10588 33746 -10574
rect 19042 -10598 33746 -10588
rect 34530 -10608 43859 -10586
rect 34530 -10700 43692 -10608
rect 43800 -10700 43859 -10608
rect 34530 -10732 43859 -10700
rect 33850 -10874 33940 -10842
rect 33850 -10942 33864 -10874
rect 33928 -10942 33940 -10874
rect 33850 -10956 33940 -10942
rect 35864 -10880 74600 -10870
rect 35864 -10942 35876 -10880
rect 35946 -10942 74450 -10880
rect 35864 -10944 74450 -10942
rect 74554 -10944 74600 -10880
rect 35864 -10955 74600 -10944
rect 34506 -11114 35694 -10968
rect 34506 -11116 34624 -11114
rect 34506 -11184 34598 -11116
rect 34506 -11248 34516 -11184
rect 34581 -11248 34598 -11184
rect 59740 -11212 59922 -11168
rect 59740 -11232 59788 -11212
rect 34506 -11264 34598 -11248
rect 35022 -11238 59788 -11232
rect 35022 -11294 35030 -11238
rect 35086 -11282 59788 -11238
rect 59884 -11282 59922 -11212
rect 35086 -11294 59922 -11282
rect 35022 -11300 59922 -11294
rect 35022 -11302 35102 -11300
rect 34730 -11344 34878 -11316
rect 59740 -11328 59922 -11300
rect 34730 -11412 34768 -11344
rect 34836 -11412 34878 -11344
rect 34730 -11452 34878 -11412
<< via3 >>
rect 5384 -9654 5518 -9522
rect 57032 -9600 57114 -9528
rect 74282 -9750 74348 -9684
rect 87118 -9930 87220 -9866
rect 1814 -10286 2230 -10092
rect 34741 -10450 34806 -10428
rect 34741 -10492 34778 -10450
rect 34778 -10492 34806 -10450
rect 19056 -10588 19120 -10524
rect 43692 -10700 43800 -10608
rect 33864 -10875 33928 -10874
rect 33864 -10941 33928 -10875
rect 33864 -10942 33928 -10941
rect 74450 -10944 74554 -10880
rect 34516 -11248 34581 -11184
rect 59788 -11282 59884 -11212
rect 34768 -11412 34836 -11344
<< metal4 >>
rect 1811 -9792 2017 133
rect 19048 -8601 19128 52
rect 5363 -9522 5550 -9500
rect 5363 -9654 5384 -9522
rect 5518 -9654 5550 -9522
rect 1762 -10092 2288 -9792
rect 1762 -10286 1814 -10092
rect 2230 -10286 2288 -10092
rect 1762 -10320 2288 -10286
rect 5363 -23086 5550 -9654
rect 19040 -10524 19130 -8601
rect 34726 -10318 34836 111
rect 34724 -10428 34836 -10318
rect 34724 -10492 34741 -10428
rect 34806 -10492 34836 -10428
rect 34724 -10514 34836 -10492
rect 19040 -10588 19056 -10524
rect 19120 -10588 19130 -10524
rect 43665 -10538 43819 99
rect 57016 11 57485 133
rect 57016 -9400 57138 11
rect 74248 -150 74398 452
rect 56994 -9462 57188 -9400
rect 56992 -9528 57188 -9462
rect 56992 -9600 57032 -9528
rect 57114 -9600 57188 -9528
rect 74280 -9556 74352 -150
rect 56992 -9644 57188 -9600
rect 56994 -9650 57188 -9644
rect 74202 -9684 74432 -9556
rect 74202 -9750 74282 -9684
rect 74348 -9750 74432 -9684
rect 74202 -9816 74432 -9750
rect 87071 -9854 87301 477
rect 87071 -9866 87300 -9854
rect 87071 -9930 87118 -9866
rect 87220 -9930 87300 -9866
rect 87071 -9938 87300 -9930
rect 19040 -10602 19130 -10588
rect 43652 -10608 43854 -10538
rect 43652 -10700 43692 -10608
rect 43800 -10700 43854 -10608
rect 43652 -10734 43854 -10700
rect 33850 -10874 33940 -10842
rect 33850 -10942 33864 -10874
rect 33928 -10942 33940 -10874
rect 33850 -10966 33940 -10942
rect 74424 -10880 74600 -10870
rect 74424 -10944 74450 -10880
rect 74554 -10944 74600 -10880
rect 74424 -10955 74600 -10944
rect 74474 -10966 74544 -10955
rect 33849 -10995 33940 -10966
rect 33849 -17566 33913 -10995
rect 5346 -23274 5550 -23086
rect 24314 -17630 33913 -17566
rect 34500 -11184 34598 -11156
rect 34500 -11248 34516 -11184
rect 34581 -11248 34598 -11184
rect 5346 -24994 5514 -23274
rect 24314 -25006 24378 -17630
rect 34500 -24943 34598 -11248
rect 59740 -11212 59926 -11186
rect 59740 -11282 59788 -11212
rect 59884 -11282 59926 -11212
rect 34732 -11344 34878 -11316
rect 59740 -11328 59926 -11282
rect 34732 -11412 34768 -11344
rect 34836 -11412 34878 -11344
rect 34732 -11452 34878 -11412
rect 34758 -17488 34842 -11452
rect 34758 -17572 43404 -17488
rect 43320 -25008 43404 -17572
rect 59795 -25033 59861 -11328
rect 74477 -25503 74544 -10966
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_11 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1611950381
transform 1 0 540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_10
timestamp 1611950381
transform 1 0 14540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_9
timestamp 1611950381
transform 1 0 28540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_8
timestamp 1611950381
transform 1 0 42540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_7
timestamp 1611950381
transform 1 0 56540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_6
timestamp 1611950381
transform 1 0 70540 0 -1 -25460
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_13
timestamp 1611950381
transform 1 0 84540 0 -1 -25460
box -540 -540 12540 14540
use sky130_fd_sc_hd__tap_1  sky130_fd_sc_hd__tap_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1611950381
transform 1 0 34106 0 -1 -9590
box -38 -48 130 592
use BITCELL  BITCELL_1
timestamp 1611860754
transform 1 0 34601 0 1 -10949
box 515 -167 1083 753
use BITCELL  BITCELL_0
timestamp 1611860754
transform 1 0 33491 0 1 -10948
box 515 -167 1083 753
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_0
timestamp 1611950381
transform 1 0 540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_1
timestamp 1611950381
transform 1 0 14540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_3
timestamp 1611950381
transform 1 0 28540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_2
timestamp 1611950381
transform 1 0 42540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_5
timestamp 1611950381
transform 1 0 56540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_4
timestamp 1611950381
transform 1 0 70540 0 1 540
box -540 -540 12540 14540
use sky130_ef_io__bare_pad  sky130_ef_io__bare_pad_12
timestamp 1611950381
transform 1 0 84540 0 1 540
box -540 -540 12540 14540
<< labels >>
flabel space 384 390 384 390 1 FreeSans 6400 0 0 0 VDD
flabel space 28406 392 28406 392 1 FreeSans 6400 0 0 0 SENSE_N
flabel space 42400 400 42400 400 1 FreeSans 6400 0 0 0 BLB
flabel space 418 -39598 418 -39598 1 FreeSans 6400 0 0 0 VSS
flabel space 28410 -39596 28410 -39596 1 FreeSans 6400 0 0 0 BL
flabel space 14394 396 14394 396 1 FreeSans 6400 0 0 0 Q0
flabel space 14398 -39602 14398 -39600 1 FreeSans 6400 0 0 0 WRR0
flabel space 42398 -39602 42398 -39602 1 FreeSans 6400 0 0 0 WRL0
flabel space 56408 402 56408 402 1 FreeSans 6400 0 0 0 Q0_N
flabel space 56400 -39598 56400 -39598 1 FreeSans 6400 0 0 0 WRR1
flabel space 70416 -39584 70416 -39584 1 FreeSans 6400 0 0 0 WRL1
flabel space 70402 400 70402 400 1 FreeSans 6400 0 0 0 Q1
flabel space 84398 402 84398 402 1 FreeSans 6400 0 0 0 Q1_N
<< end >>
