magic
tech sky130A
magscale 1 2
timestamp 1612374967
<< nmos >>
rect 652 -139 682 -19
rect 740 -139 770 -19
rect 828 -139 858 -19
rect 916 -139 946 -19
<< ndiff >>
rect 594 -60 652 -19
rect 594 -94 606 -60
rect 640 -94 652 -60
rect 594 -139 652 -94
rect 682 -60 740 -19
rect 682 -94 694 -60
rect 728 -94 740 -60
rect 682 -139 740 -94
rect 770 -60 828 -19
rect 770 -94 782 -60
rect 816 -94 828 -60
rect 770 -139 828 -94
rect 858 -60 916 -19
rect 858 -94 870 -60
rect 904 -94 916 -60
rect 858 -139 916 -94
rect 946 -60 1004 -19
rect 946 -94 958 -60
rect 992 -94 1004 -60
rect 946 -139 1004 -94
<< ndiffc >>
rect 606 -94 640 -60
rect 694 -94 728 -60
rect 782 -94 816 -60
rect 870 -94 904 -60
rect 958 -94 992 -60
<< poly >>
rect 515 46 581 63
rect 515 12 531 46
rect 565 35 581 46
rect 1015 47 1081 64
rect 1015 35 1031 47
rect 565 12 770 35
rect 515 -3 770 12
rect 515 -4 581 -3
rect 652 -19 682 -3
rect 740 -19 770 -3
rect 828 13 1031 35
rect 1065 13 1081 47
rect 828 -3 1081 13
rect 828 -19 858 -3
rect 916 -19 946 -3
rect 652 -165 682 -139
rect 740 -165 770 -139
rect 828 -165 858 -139
rect 916 -165 946 -139
<< polycont >>
rect 531 12 565 46
rect 1031 13 1065 47
<< locali >>
rect 694 113 728 123
rect 708 97 728 113
rect 871 97 904 125
rect 531 46 565 63
rect 531 -5 565 12
rect 606 -60 640 -19
rect 606 -129 640 -102
rect 694 -60 728 97
rect 694 -128 728 -102
rect 782 -60 816 -19
rect 782 -128 816 -102
rect 870 -60 904 97
rect 1031 47 1065 64
rect 1031 -4 1065 13
rect 870 -128 904 -102
rect 958 -60 992 -19
rect 958 -128 992 -102
<< viali >>
rect 606 -94 640 -68
rect 606 -102 640 -94
rect 694 -94 728 -68
rect 694 -102 728 -94
rect 782 -94 816 -68
rect 782 -102 816 -94
rect 870 -94 904 -68
rect 870 -102 904 -94
rect 958 -94 992 -68
rect 958 -102 992 -94
<< metal1 >>
rect 676 87 746 95
rect 676 35 684 87
rect 736 35 746 87
rect 676 29 746 35
rect 853 87 923 95
rect 853 35 864 87
rect 916 35 923 87
rect 853 29 923 35
rect 594 -59 647 -19
rect 646 -111 647 -59
rect 594 -139 647 -111
rect 682 -68 740 29
rect 682 -102 694 -68
rect 728 -102 740 -68
rect 682 -140 740 -102
rect 772 -59 825 -19
rect 824 -111 825 -59
rect 772 -139 825 -111
rect 858 -68 916 29
rect 858 -102 870 -68
rect 904 -102 916 -68
rect 858 -140 916 -102
rect 951 -59 1004 -19
rect 1003 -111 1004 -59
rect 951 -139 1004 -111
<< via1 >>
rect 684 35 736 87
rect 864 35 916 87
rect 594 -68 646 -59
rect 594 -102 606 -68
rect 606 -102 640 -68
rect 640 -102 646 -68
rect 594 -111 646 -102
rect 772 -68 824 -59
rect 772 -102 782 -68
rect 782 -102 816 -68
rect 816 -102 824 -68
rect 772 -111 824 -102
rect 951 -68 1003 -59
rect 951 -102 958 -68
rect 958 -102 992 -68
rect 992 -102 1003 -68
rect 951 -111 1003 -102
<< metal2 >>
rect 677 126 771 155
rect 677 95 695 126
rect 676 87 695 95
rect 676 35 684 87
rect 751 70 771 126
rect 736 35 771 70
rect 676 29 771 35
rect 677 28 771 29
rect 828 126 922 154
rect 828 70 849 126
rect 905 96 922 126
rect 905 87 923 96
rect 828 35 864 70
rect 916 35 923 87
rect 828 29 923 35
rect 828 27 922 29
rect 594 -57 659 -19
rect 650 -113 659 -57
rect 594 -139 659 -113
rect 762 -57 835 -19
rect 762 -113 771 -57
rect 827 -113 835 -57
rect 762 -139 835 -113
rect 941 -57 1004 -19
rect 941 -113 948 -57
rect 941 -139 1004 -113
<< via2 >>
rect 695 87 751 126
rect 695 70 736 87
rect 736 70 751 87
rect 849 87 905 126
rect 849 70 864 87
rect 864 70 905 87
rect 594 -59 650 -57
rect 594 -111 646 -59
rect 646 -111 650 -59
rect 594 -113 650 -111
rect 771 -59 827 -57
rect 771 -111 772 -59
rect 772 -111 824 -59
rect 824 -111 827 -59
rect 771 -113 827 -111
rect 948 -59 1004 -57
rect 948 -111 951 -59
rect 951 -111 1003 -59
rect 1003 -111 1004 -59
rect 948 -113 1004 -111
<< metal3 >>
rect 532 317 1077 364
rect 532 253 692 317
rect 756 253 843 317
rect 907 253 1077 317
rect 532 214 1077 253
rect 676 126 768 154
rect 676 70 695 126
rect 751 70 768 126
rect 676 43 768 70
rect 831 126 924 154
rect 831 70 849 126
rect 905 70 924 126
rect 831 41 924 70
rect 573 -57 1083 -19
rect 573 -113 594 -57
rect 650 -113 771 -57
rect 827 -113 948 -57
rect 1004 -113 1083 -57
rect 573 -167 1083 -113
<< via3 >>
rect 692 253 756 317
rect 843 253 907 317
<< metal4 >>
rect 680 317 768 348
rect 680 253 692 317
rect 756 253 768 317
rect 680 42 768 253
rect 832 317 920 348
rect 832 253 843 317
rect 907 253 920 317
rect 832 42 920 253
use SENSEAMP  SENSEAMP_0
timestamp 1612374967
transform 1 0 558 0 1 459
box 0 -370 482 294
<< end >>
