magic
tech sky130A
magscale 1 2
timestamp 1611715700
<< nwell >>
rect -109 -117 109 117
<< pmos >>
rect -15 -55 15 55
<< pdiff >>
rect -73 43 -15 55
rect -73 -43 -61 43
rect -27 -43 -15 43
rect -73 -55 -15 -43
rect 15 43 73 55
rect 15 -43 27 43
rect 61 -43 73 43
rect 15 -55 73 -43
<< pdiffc >>
rect -61 -43 -27 43
rect 27 -43 61 43
<< poly >>
rect -15 55 15 81
rect -15 -81 15 -55
<< locali >>
rect -61 43 -27 59
rect -61 -59 -27 -43
rect 27 43 61 59
rect 27 -59 61 -43
<< viali >>
rect -61 -43 -27 43
rect 27 -43 61 43
<< metal1 >>
rect -67 43 -21 55
rect -67 -43 -61 43
rect -27 -43 -21 43
rect -67 -55 -21 -43
rect 21 43 67 55
rect 21 -43 27 43
rect 61 -43 67 43
rect 21 -55 67 -43
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 0.55 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
