magic
tech sky130A
magscale 1 2
timestamp 1611776490
<< nmos >>
rect -120 -60 -90 60
rect 90 -60 120 60
<< ndiff >>
rect -178 29 -120 60
rect -182 17 -120 29
rect -182 -17 -170 17
rect -136 -17 -120 17
rect -182 -29 -120 -17
rect -178 -60 -120 -29
rect -90 29 -32 60
rect 32 29 90 60
rect -90 17 -28 29
rect -90 -17 -74 17
rect -40 -17 -28 17
rect -90 -29 -28 -17
rect 28 17 90 29
rect 28 -17 40 17
rect 74 -17 90 17
rect 28 -29 90 -17
rect -90 -60 -32 -29
rect 32 -60 90 -29
rect 120 29 178 60
rect 120 17 182 29
rect 120 -17 136 17
rect 170 -17 182 17
rect 120 -29 182 -17
rect 120 -60 178 -29
<< ndiffc >>
rect -170 -17 -136 17
rect -74 -17 -40 17
rect 40 -17 74 17
rect 136 -17 170 17
<< poly >>
rect 72 132 138 148
rect 72 98 88 132
rect 122 98 138 132
rect -120 60 -90 86
rect 72 82 138 98
rect 90 60 120 82
rect -120 -82 -90 -60
rect -138 -98 -72 -82
rect 90 -86 120 -60
rect -138 -132 -122 -98
rect -88 -132 -72 -98
rect -138 -148 -72 -132
<< polycont >>
rect 88 98 122 132
rect -122 -132 -88 -98
<< locali >>
rect 72 98 88 132
rect 122 98 138 132
rect -170 17 -136 33
rect -170 -33 -136 -17
rect -74 17 -40 33
rect -74 -33 -40 -17
rect 40 17 74 33
rect 40 -33 74 -17
rect 136 17 170 33
rect 136 -33 170 -17
rect -138 -132 -122 -98
rect -88 -132 -72 -98
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 0.6 l 0.150 m 1 nf 2 diffcov 20 polycov 20 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 0 rlcov 0 topc 0 botc 0 poverlap 1 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt} full_metal 0 viasrc 0 viadrn 0 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
