magic
tech sky130A
magscale 1 2
timestamp 1611860754
<< nmos >>
rect 652 -139 682 -19
rect 740 -139 770 -19
rect 828 -139 858 -19
rect 916 -139 946 -19
<< ndiff >>
rect 594 -42 652 -19
rect 594 -112 606 -42
rect 640 -112 652 -42
rect 594 -139 652 -112
rect 682 -42 740 -19
rect 682 -112 694 -42
rect 728 -112 740 -42
rect 682 -139 740 -112
rect 770 -42 828 -19
rect 770 -112 782 -42
rect 816 -112 828 -42
rect 770 -139 828 -112
rect 858 -42 916 -19
rect 858 -112 870 -42
rect 904 -112 916 -42
rect 858 -139 916 -112
rect 946 -42 1004 -19
rect 946 -112 958 -42
rect 992 -112 1004 -42
rect 946 -139 1004 -112
<< ndiffc >>
rect 606 -112 640 -42
rect 694 -112 728 -42
rect 782 -112 816 -42
rect 870 -112 904 -42
rect 958 -112 992 -42
<< poly >>
rect 515 46 581 63
rect 515 12 531 46
rect 565 35 581 46
rect 1015 47 1081 64
rect 1015 35 1031 47
rect 565 12 770 35
rect 515 -3 770 12
rect 515 -4 581 -3
rect 652 -19 682 -3
rect 740 -19 770 -3
rect 828 13 1031 35
rect 1065 13 1081 47
rect 828 -3 1081 13
rect 828 -19 858 -3
rect 916 -19 946 -3
rect 652 -165 682 -139
rect 740 -165 770 -139
rect 828 -165 858 -139
rect 916 -165 946 -139
<< polycont >>
rect 531 12 565 46
rect 1031 13 1065 47
<< locali >>
rect 694 113 728 123
rect 708 97 728 113
rect 871 97 904 125
rect 531 46 565 63
rect 531 -5 565 12
rect 606 -42 640 -19
rect 606 -129 640 -127
rect 694 -42 728 97
rect 694 -128 728 -127
rect 782 -42 816 -19
rect 782 -128 816 -127
rect 870 -42 904 97
rect 1031 47 1065 64
rect 1031 -4 1065 13
rect 870 -128 904 -127
rect 958 -42 992 -19
rect 958 -128 992 -127
<< viali >>
rect 606 -112 640 -42
rect 606 -127 640 -112
rect 694 -112 728 -42
rect 694 -127 728 -112
rect 782 -112 816 -42
rect 782 -127 816 -112
rect 870 -112 904 -42
rect 870 -127 904 -112
rect 958 -112 992 -42
rect 958 -127 992 -112
<< metal1 >>
rect 676 87 746 95
rect 676 35 684 87
rect 736 35 746 87
rect 676 29 746 35
rect 853 89 923 95
rect 853 34 864 89
rect 916 34 923 89
rect 853 29 923 34
rect 594 -42 647 -19
rect 594 -139 647 -127
rect 682 -42 740 29
rect 682 -127 694 -42
rect 728 -127 740 -42
rect 682 -140 740 -127
rect 772 -42 825 -19
rect 772 -139 825 -127
rect 858 -42 916 29
rect 858 -127 870 -42
rect 904 -127 916 -42
rect 858 -140 916 -127
rect 951 -42 1004 -19
rect 951 -139 1004 -127
<< via1 >>
rect 684 35 736 87
rect 864 34 916 89
rect 594 -127 606 -42
rect 606 -127 640 -42
rect 640 -127 647 -42
rect 772 -127 782 -42
rect 782 -127 816 -42
rect 816 -127 825 -42
rect 951 -127 958 -42
rect 958 -127 992 -42
rect 992 -127 1004 -42
<< metal2 >>
rect 677 145 771 155
rect 677 95 687 145
rect 676 87 687 95
rect 676 35 684 87
rect 759 52 771 145
rect 736 35 771 52
rect 676 29 771 35
rect 677 28 771 29
rect 828 145 922 154
rect 828 52 841 145
rect 913 96 922 145
rect 913 89 923 96
rect 828 34 864 52
rect 916 34 923 89
rect 828 29 923 34
rect 828 27 922 29
rect 594 -42 659 -19
rect 650 -128 659 -42
rect 594 -139 659 -128
rect 762 -42 835 -19
rect 762 -128 771 -42
rect 827 -128 835 -42
rect 762 -139 835 -128
rect 941 -42 1004 -19
rect 941 -127 948 -42
rect 941 -139 1004 -127
<< via2 >>
rect 687 87 759 145
rect 687 52 736 87
rect 736 52 759 87
rect 841 89 913 145
rect 841 52 864 89
rect 864 52 913 89
rect 594 -127 647 -42
rect 647 -127 650 -42
rect 594 -128 650 -127
rect 771 -127 772 -42
rect 772 -127 825 -42
rect 825 -127 827 -42
rect 771 -128 827 -127
rect 948 -127 951 -42
rect 951 -127 1004 -42
<< metal3 >>
rect 532 338 1077 364
rect 532 233 692 338
rect 757 233 843 338
rect 908 233 1077 338
rect 532 214 1077 233
rect 676 145 768 154
rect 676 52 687 145
rect 759 52 768 145
rect 676 43 768 52
rect 831 145 924 154
rect 831 52 841 145
rect 913 52 924 145
rect 831 41 924 52
rect 573 -42 1083 -19
rect 573 -128 594 -42
rect 650 -128 771 -42
rect 827 -127 948 -42
rect 1004 -127 1083 -42
rect 827 -128 1083 -127
rect 573 -167 1083 -128
<< via3 >>
rect 692 233 757 338
rect 843 233 908 338
<< mtj >>
rect 708 93 728 113
rect 870 93 890 113
<< metal4 >>
rect 680 338 768 348
rect 680 233 692 338
rect 757 233 768 338
rect 680 42 768 233
rect 832 338 920 348
rect 832 233 843 338
rect 908 233 920 338
rect 832 42 920 233
use SENSEAMP  SENSEAMP_0
timestamp 1611851455
transform 1 0 558 0 1 459
box 0 -370 482 294
<< end >>
